CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 15 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
11
7 Pulser~
4 110 335 0 10 12
0 27 28 15 29 0 0 5 5 1
8
0
0 0 4640 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3780 0 0
2
43530.4 10
0
2 +V
167 171 147 0 1 3
0 17
0
0 0 54240 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9265 0 0
2
43530.4 9
0
6 74LS48
188 888 257 0 14 29
0 9 10 11 12 24 25 2 3 4
5 6 7 8 26
0
0 0 4832 0
7 74LS248
-24 -60 25 -52
2 U4
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9442 0 0
2
43530.4 8
0
6 74112~
219 329 253 0 7 32
0 17 16 15 16 17 23 12
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 3 0
1 U
9424 0 0
2
43530.4 7
0
6 74112~
219 435 253 0 7 32
0 17 12 15 12 17 22 11
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 3 0
1 U
9968 0 0
2
43530.4 6
0
6 74112~
219 544 248 0 7 32
0 17 14 15 14 17 21 10
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
9281 0 0
2
43530.4 5
0
6 74112~
219 644 247 0 7 32
0 17 13 15 13 17 20 9
0
0 0 4704 0
5 74112
4 -60 39 -52
3 U2A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
8464 0 0
2
43530.4 4
0
9 2-In AND~
219 430 74 0 3 22
0 12 11 14
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7168 0 0
2
43530.4 3
0
9 2-In AND~
219 580 75 0 3 22
0 14 10 13
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3171 0 0
2
43530.4 2
0
9 CC 7-Seg~
183 1063 225 0 18 19
10 8 7 6 5 4 3 2 18 19
0 0 0 0 0 0 0 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
4139 0 0
2
43530.4 1
0
13 Logic Switch~
5 148 211 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6435 0 0
2
43530.4 0
0
37
7 7 2 0 0 0 0 3 10 0 0 5
920 221
1013 221
1013 294
1078 294
1078 261
8 6 3 0 0 0 0 3 10 0 0 5
920 230
1018 230
1018 289
1072 289
1072 261
9 5 4 0 0 0 0 3 10 0 0 5
920 239
1023 239
1023 284
1066 284
1066 261
10 4 5 0 0 0 0 3 10 0 0 5
920 248
1028 248
1028 279
1060 279
1060 261
11 3 6 0 0 0 0 3 10 0 0 5
920 257
1033 257
1033 269
1054 269
1054 261
12 2 7 0 0 0 0 3 10 0 0 3
920 266
1048 266
1048 261
13 1 8 0 0 0 0 3 10 0 0 3
920 275
1042 275
1042 261
7 1 9 0 0 0 0 7 3 0 0 4
668 211
843 211
843 221
856 221
0 2 10 0 0 0 0 0 3 14 0 6
579 206
600 206
600 269
838 269
838 230
856 230
0 3 11 0 0 0 0 0 3 18 0 4
473 265
843 265
843 239
856 239
7 4 12 0 0 0 0 4 3 0 0 6
353 217
367 217
367 177
848 177
848 248
856 248
0 4 13 0 0 0 0 0 7 13 0 3
606 117
606 229
620 229
3 2 13 0 0 0 0 9 7 0 0 4
601 75
606 75
606 211
620 211
2 7 10 0 0 0 0 9 6 0 0 6
556 84
552 84
552 181
579 181
579 212
568 212
0 4 14 0 0 0 0 0 6 17 0 3
469 74
469 230
520 230
0 1 14 0 0 0 0 0 9 17 0 3
505 74
505 66
556 66
3 2 14 0 0 0 0 8 6 0 0 4
451 74
506 74
506 212
520 212
2 7 11 0 0 0 0 8 5 0 0 6
406 83
396 83
396 270
473 270
473 217
459 217
1 0 12 0 0 0 0 8 0 0 25 3
406 65
375 65
375 217
3 0 15 0 0 0 0 7 0 0 23 3
614 220
610 220
610 326
3 0 15 0 0 0 0 6 0 0 23 3
514 221
510 221
510 326
3 0 15 0 0 0 0 5 0 0 23 3
405 226
401 226
401 326
0 0 15 0 0 0 0 0 0 26 0 2
291 326
730 326
0 4 12 0 0 0 0 0 5 25 0 3
383 217
383 235
411 235
0 2 12 0 0 0 0 0 5 0 0 2
366 217
411 217
3 3 15 0 0 0 0 1 4 0 0 4
134 326
291 326
291 226
299 226
0 4 16 0 0 0 0 0 4 28 0 3
184 217
184 235
305 235
1 2 16 0 0 16 0 11 4 0 0 3
160 211
160 217
305 217
5 0 17 0 0 0 0 4 0 0 37 2
329 265
329 296
5 0 17 0 0 0 0 7 0 0 37 2
644 259
644 296
5 0 17 0 0 0 0 6 0 0 37 2
544 260
544 296
5 0 17 0 0 0 0 5 0 0 37 2
435 265
435 296
0 1 17 0 0 0 0 0 7 37 0 2
644 156
644 184
0 1 17 0 0 0 0 0 6 37 0 2
544 156
544 185
1 0 17 0 0 0 0 5 0 0 37 2
435 190
435 156
0 1 17 0 0 0 0 0 4 37 0 3
327 156
329 156
329 190
1 0 17 0 0 0 0 2 0 0 0 4
171 156
731 156
731 296
171 296
1
-16 0 0 0 400 0 0 0 0 3 2 1 18
8 Elephant
0 0 0 24
208 360 422 391
219 368 410 389
24 Gudito, Steaven Klein F.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
